begin

J1 <= Q2 AND X;
K1 <= (NOT Q2) OR X;
J2 <= X;
K2 <= NOT X;
Z <= Q1 AND (NOT Q2) AND X;

end Behavioral;
